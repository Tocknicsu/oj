module tb;
reg CLK, RESET, ADD, SUB;
